module decode(
    input wire clk,
    input wire rst,
    input wire[31:0] instr
);


endmodule