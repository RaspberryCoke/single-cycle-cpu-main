module execute(
    input wire clk,
    input wire rst,
    input wire[31:0] instr
);


endmodule

